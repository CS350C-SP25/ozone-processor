import uop_pkg::*;
import reg_pkg::*;
import is_pkg::*;

