// used for the RAT + RRAT