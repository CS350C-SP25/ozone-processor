module branch_pred #(
    //gay sex
) (
    //more gay sex
);
    //epic amounts of gay sex
endmodule