package reg_pkg;
    parameter int NUM_ARCH_REGS = 32; // x0-x31 as per RISC-V
    parameter int ADDR_BITS = 64;
endpackage