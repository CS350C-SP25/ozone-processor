import uop_pkg::*;
import reg_pkg::*;
import ins_sched_pkg::*;

