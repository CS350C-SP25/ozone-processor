module #(
    
) backend();

endmodule: backend