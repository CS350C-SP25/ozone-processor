`ifndef MEM_PKG_SV
`define MEM_PKG_SV
package mem_pkg;
  parameter int LQ_SIZE = 32;
endpackage
`endif // MEM_PKG_SV
