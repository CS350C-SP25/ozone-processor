`include "./"
module #(
    
) backend();

endmodule: backend